** test dac 3 bits

.include tsmc_spice_model.txt
.include inverter.cir
.include dac_3.cir

Vdd vdd gnd 1.8V//PULSE(1.8 0 0 0.1n 0.1n 2.5n 5n)
*Vin in gnd SIN(0.9 0.9 20MEG 0 0)
*Vdummy 1 gnd 0V
*V0 out0 gnd 0
*V1 out1 gnd 0
*V2 out2 gnd 0

************ lsb  1  msb**********
xdac vdd gnd vdd vdd vdd out dac_3


.control
save all @xadc.Mn_sw1_1[id]
tran 1n 50n
.endc
.END